----------------------------------------------------------------------------------
-- Ecole : 					INSA Toulouse
-- Etudiants : 			Laure FEUILLET et Maël PLANTEC
--
-- Nom du projet :	Projet Système Informatique
-- Module :	        Test de la pipeline
----------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY test_pipeline IS
END test_pipeline;

ARCHITECTURE behavior OF test_pipeline IS
    -- Component Declaration for the Unit Under Test (UUT)
    COMPONENT Pipeline
    PORT(
         Ck : IN  std_logic;
         OPi : IN  std_logic_vector(7 downto 0);
         Ai : IN  std_logic_vector(15 downto 0);
         Bi : IN  std_logic_vector(15 downto 0);
         Ci : IN  std_logic_vector(15 downto 0);
         OPo : OUT  std_logic_vector(7 downto 0);
         Ao : OUT  std_logic_vector(15 downto 0);
         Bo : OUT  std_logic_vector(15 downto 0);
         Co : OUT  std_logic_vector(15 downto 0)
        );
    END COMPONENT;

   --Inputs
   signal Ck : std_logic := '0';
   signal OPi : std_logic_vector(7 downto 0) := (others => '0');
   signal Ai : std_logic_vector(15 downto 0) := (others => '0');
   signal Bi : std_logic_vector(15 downto 0) := (others => '0');
   signal Ci : std_logic_vector(15 downto 0) := (others => '0');
 	--Outputs
   signal OPo : std_logic_vector(7 downto 0);
   signal Ao : std_logic_vector(15 downto 0);
   signal Bo : std_logic_vector(15 downto 0);
   signal Co : std_logic_vector(15 downto 0);
   -- Clock
   constant Ck_period : time := 10 ns;

BEGIN
	-- Instantiate the Unit Under Test (UUT)
   uut: Pipeline PORT MAP (
          Ck => Ck,
          OPi => OPi,
          Ai => Ai,
          Bi => Bi,
          Ci => Ci,
          OPo => OPo,
          Ao => Ao,
          Bo => Bo,
          Co => Co
        );
   -- Clock process definitions
   Ck_process :process
   begin
		Ck <= '0';
		wait for Ck_period/2;
		Ck <= '1';
		wait for Ck_period/2;
   end process;

   -- Stimulus process
   stim_proc: process
   begin
    wait for 100 ns;
		OPi <= x"01";
		Ai <= x"0002";
		Bi <= x"0003";
		Ci <= x"0004";

    wait;
   end process;
END;
